module happy(SW,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7); 
input [3:0]SW; 
output reg[6:0]HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7; 
always @ (SW) 
begin 
case (SW) 
4'b0000: begin 
HEX7 =7'b 0010001; //Y
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
end 
4'b0001: begin 
HEX7 =7'b 0001100; //P
HEX6 =7'b 0010001; //Y
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
 end 
4'b0010: begin 
HEX7 =7'b 0001100; //P
HEX6 =7'b 0001100; //P
HEX5 =7'b 0010001; //Y
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
end 
4'b0011: begin 
HEX7 =7'b 0001000; //A
HEX6 =7'b 0001100; //P
HEX5 =7'b 0001100; //P
HEX4 =7'b 0010001; //Y
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
end 
4'b0100: begin 
HEX7 =7'b 0001001; //H
HEX6 =7'b 0001000; //A
HEX5 =7'b 0001100; //P
HEX4 =7'b 0001100; //P
HEX3 =7'b 0010001; //Y
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
end 
4'b0101: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 0001001; //H
HEX5 =7'b 0001000; //A
HEX4 =7'b 0001100; //P
HEX3 =7'b 0001100; //P
HEX2 =7'b 0010001; //Y
HEX1 =7'b 1111111;
HEX0 =7'b 1111111;
end 
4'b0110: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 0001001; //H
HEX4 =7'b 0001000; //A
HEX3 =7'b 0001100; //P
HEX2 =7'b 0001100; //P
HEX1 =7'b 0010001; //Y
HEX0 =7'b 1111111; 
end 
4'b0111: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 0001001; //H
HEX3 =7'b 0001000; //A
HEX2 =7'b 0001100; //P
HEX1 =7'b 0001100; //P
HEX0 =7'b 0010001; //Y
end 
4'b1000: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 0001001; //H
HEX2 =7'b 0001000; //A
HEX1 =7'b 0001100; //P
HEX0 =7'b 0001100; //P
end 
4'b1001: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 0001001; //H
HEX1 =7'b 0001000; //A
HEX0 =7'b 0001100; //P
end 
4'b1010: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 0001001; //H
HEX0 =7'b 0001000; //A
end 
4'b1011: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 0001001; //H
end 
4'b1100: begin 
HEX7 =7'b 1111111;
HEX6 =7'b 1111111;
HEX5 =7'b 1111111;
HEX4 =7'b 1111111;
HEX3 =7'b 1111111;
HEX2 =7'b 1111111;
HEX1 =7'b 1111111;
HEX0 =7'b 1111111; 
end 
endcase 
end 
endmodule 